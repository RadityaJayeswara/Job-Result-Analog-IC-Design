magic
tech sky130A
magscale 1 2
timestamp 1729394227
<< nwell >>
rect 1494 1521 3258 1768
rect 1494 1498 2203 1521
rect 2253 1515 3258 1521
rect 2253 1498 2499 1515
rect 1494 1496 2499 1498
rect 2533 1496 3258 1515
rect 1494 1400 3258 1496
rect 1494 1364 1908 1400
rect 1962 1364 3258 1400
rect 1494 1274 3258 1364
rect 1494 1249 2207 1274
rect 2252 1249 3258 1274
rect 1494 1033 3258 1249
rect 1494 998 1912 1033
rect 1971 1030 3258 1033
rect 1971 1008 2206 1030
rect 2252 1008 2494 1030
rect 1971 1003 2494 1008
rect 2547 1003 3258 1030
rect 1971 998 3258 1003
rect 1494 938 3258 998
rect 1494 906 1912 938
rect 1954 926 3258 938
rect 1954 914 2774 926
rect 2806 914 3258 926
rect 1954 906 2766 914
rect 1494 854 2766 906
rect 2830 854 3258 914
rect 1494 509 3258 854
<< nsubdiff >>
rect 1530 1698 1590 1732
rect 3162 1698 3222 1732
rect 1530 1672 1564 1698
rect 3188 1672 3222 1698
rect 1530 579 1564 605
rect 3188 579 3222 605
rect 1530 545 1590 579
rect 3162 545 3222 579
<< nsubdiffcont >>
rect 1590 1698 3162 1732
rect 1530 605 1564 1672
rect 3188 605 3222 1672
rect 1590 545 3162 579
<< poly >>
rect 1614 1564 1706 1580
rect 1614 1530 1630 1564
rect 1664 1530 1706 1564
rect 1614 1514 1706 1530
rect 1676 1509 1706 1514
rect 3046 1564 3138 1580
rect 3046 1530 3088 1564
rect 3122 1530 3138 1564
rect 3046 1514 3138 1530
rect 3046 1509 3076 1514
rect 1676 765 1706 770
rect 1614 749 1706 765
rect 1614 715 1630 749
rect 1664 715 1706 749
rect 1614 699 1706 715
rect 3046 765 3076 770
rect 3046 749 3138 765
rect 3046 715 3088 749
rect 3122 715 3138 749
rect 3046 699 3138 715
<< polycont >>
rect 1630 1530 1664 1564
rect 3088 1530 3122 1564
rect 1630 715 1664 749
rect 3088 715 3122 749
<< locali >>
rect 1530 1698 1590 1732
rect 3162 1698 3222 1732
rect 1530 1672 1564 1698
rect 3188 1672 3222 1698
rect 1614 1530 1630 1564
rect 1664 1530 1680 1564
rect 3072 1530 3088 1564
rect 3122 1530 3138 1564
rect 1614 715 1630 749
rect 1664 715 1680 749
rect 3072 715 3088 749
rect 3122 715 3138 749
rect 1530 579 1564 605
rect 3188 579 3222 605
rect 1530 545 1590 579
rect 3162 545 3222 579
<< viali >>
rect 2341 1630 2409 1664
rect 1630 1530 1664 1564
rect 3088 1530 3122 1564
rect 1630 715 1664 749
rect 3088 715 3122 749
rect 2342 613 2410 647
<< metal1 >>
rect 2329 1673 2421 1685
rect 2329 1621 2341 1673
rect 2409 1621 2421 1673
rect 2329 1573 2421 1621
rect 1618 1564 1676 1570
rect 1618 1530 1630 1564
rect 1664 1530 1676 1564
rect 1618 1524 1676 1530
rect 1630 1483 1664 1524
rect 1900 1521 1910 1573
rect 1978 1521 1988 1573
rect 2194 1521 2558 1573
rect 2764 1521 2774 1573
rect 2842 1521 2852 1573
rect 3076 1564 3134 1570
rect 3076 1530 3088 1564
rect 3122 1530 3134 1564
rect 3076 1524 3134 1530
rect 3088 1483 3122 1524
rect 1630 1471 1894 1483
rect 1630 1295 1774 1471
rect 1826 1295 1894 1471
rect 1630 1283 1894 1295
rect 2000 1283 2176 1483
rect 2288 1471 2464 1483
rect 2288 1295 2350 1471
rect 2402 1295 2464 1471
rect 2288 1283 2464 1295
rect 2576 1283 2752 1483
rect 2864 1471 3128 1483
rect 2864 1295 2926 1471
rect 2978 1295 3128 1471
rect 2864 1283 3128 1295
rect 2065 1163 2111 1283
rect 2641 1163 2687 1283
rect 2065 1116 2687 1163
rect 2065 996 2111 1116
rect 2641 996 2687 1116
rect 1624 984 1888 996
rect 1624 808 1774 984
rect 1826 808 1888 984
rect 1624 796 1888 808
rect 2000 796 2176 996
rect 2288 984 2464 996
rect 2288 808 2350 984
rect 2402 808 2464 984
rect 2288 796 2464 808
rect 2576 796 2752 996
rect 2864 984 3128 996
rect 2864 808 2926 984
rect 2978 808 3128 984
rect 2864 796 3128 808
rect 1630 755 1664 796
rect 1618 749 1676 755
rect 1618 715 1630 749
rect 1664 715 1676 749
rect 1618 709 1676 715
rect 1900 706 1910 758
rect 1978 706 1988 758
rect 2194 706 2558 758
rect 2764 706 2774 758
rect 2842 706 2852 758
rect 3088 755 3122 796
rect 3076 749 3134 755
rect 3076 715 3088 749
rect 3122 715 3134 749
rect 3076 709 3134 715
rect 2330 656 2422 706
rect 2330 604 2342 656
rect 2410 604 2422 656
rect 2330 591 2422 604
<< via1 >>
rect 2341 1664 2409 1673
rect 2341 1630 2409 1664
rect 2341 1621 2409 1630
rect 1910 1521 1978 1573
rect 2774 1521 2842 1573
rect 1774 1295 1826 1471
rect 2350 1295 2402 1471
rect 2926 1295 2978 1471
rect 1774 808 1826 984
rect 2350 808 2402 984
rect 2926 808 2978 984
rect 1910 706 1978 758
rect 2774 706 2842 758
rect 2342 647 2410 656
rect 2342 613 2410 647
rect 2342 604 2410 613
<< metal2 >>
rect 2341 1675 2409 1685
rect 1613 1605 1978 1673
rect 2341 1609 2409 1619
rect 1613 666 1681 1605
rect 1910 1573 1978 1605
rect 1910 1511 1978 1521
rect 2774 1605 3139 1673
rect 2774 1573 2842 1605
rect 2774 1511 2842 1521
rect 1774 1471 1826 1481
rect 1774 1165 1826 1295
rect 2348 1471 2404 1481
rect 2348 1285 2404 1295
rect 2926 1471 2978 1481
rect 2926 1166 2978 1295
rect 2896 1165 2978 1166
rect 1774 1114 2978 1165
rect 1772 984 1828 994
rect 1772 798 1828 808
rect 2350 984 2402 1114
rect 2350 798 2402 808
rect 2924 984 2980 994
rect 2924 798 2980 808
rect 1910 760 1978 770
rect 1910 694 1978 704
rect 2774 760 2842 770
rect 2774 694 2842 704
rect 2342 666 2410 667
rect 3071 666 3139 1605
rect 1613 656 3139 666
rect 1613 604 2342 656
rect 2410 604 3139 656
rect 1613 594 3139 604
rect 2342 591 2410 594
<< via2 >>
rect 2341 1673 2409 1675
rect 2341 1621 2409 1673
rect 2341 1619 2409 1621
rect 2348 1295 2350 1471
rect 2350 1295 2402 1471
rect 2402 1295 2404 1471
rect 1772 808 1774 984
rect 1774 808 1826 984
rect 1826 808 1828 984
rect 2924 808 2926 984
rect 2926 808 2978 984
rect 2978 808 2980 984
rect 1910 758 1978 760
rect 1910 706 1978 758
rect 1910 704 1978 706
rect 2774 758 2842 760
rect 2774 706 2842 758
rect 2774 704 2842 706
<< metal3 >>
rect 1613 1675 3139 1680
rect 1613 1619 2341 1675
rect 2409 1619 3139 1675
rect 1613 1612 3139 1619
rect 1613 675 1681 1612
rect 2338 1471 2414 1476
rect 2338 1295 2348 1471
rect 2404 1295 2414 1471
rect 2338 1177 2414 1295
rect 1762 1102 2990 1177
rect 1762 984 1838 1102
rect 1762 808 1772 984
rect 1828 808 1838 984
rect 1762 803 1838 808
rect 2914 984 2990 1102
rect 2914 808 2924 984
rect 2980 808 2990 984
rect 2914 803 2990 808
rect 1900 760 1988 765
rect 1900 704 1910 760
rect 1978 704 1988 760
rect 1900 675 1988 704
rect 1613 608 1988 675
rect 2764 760 2852 765
rect 2764 704 2774 760
rect 2842 704 2852 760
rect 2764 675 2852 704
rect 3071 675 3139 1612
rect 2764 608 3139 675
use sky130_fd_pr__pfet_01v8_QKGXH2  sky130_fd_pr__pfet_01v8_QKGXH2_0
timestamp 1729233515
transform 1 0 3061 0 1 1383
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_QKGXH2  sky130_fd_pr__pfet_01v8_QKGXH2_3
timestamp 1729233515
transform 1 0 3061 0 1 896
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_QKGXH2  sky130_fd_pr__pfet_01v8_QKGXH2_4
timestamp 1729233515
transform 1 0 1691 0 1 1383
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_QKGXH2  sky130_fd_pr__pfet_01v8_QKGXH2_5
timestamp 1729233515
transform 1 0 1691 0 1 896
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_0
timestamp 1729240055
transform 1 0 2808 0 1 896
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_1
timestamp 1729240055
transform 1 0 1944 0 1 1383
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_2
timestamp 1729240055
transform 1 0 2232 0 1 1383
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_3
timestamp 1729240055
transform 1 0 2520 0 1 1383
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_4
timestamp 1729240055
transform 1 0 2808 0 1 1383
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_5
timestamp 1729240055
transform 1 0 1944 0 1 896
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_6
timestamp 1729240055
transform 1 0 2232 0 1 896
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_7
timestamp 1729240055
transform 1 0 2520 0 1 896
box -144 -200 144 200
<< labels >>
flabel metal3 1802 1028 1802 1028 0 FreeSans 160 0 0 0 D7
port 2 nsew
flabel metal2 1796 1248 1796 1248 0 FreeSans 160 0 0 0 D6
port 3 nsew
flabel metal1 2092 1238 2092 1238 0 FreeSans 160 0 0 0 D5
port 4 nsew
flabel locali 3206 1700 3206 1700 0 FreeSans 160 0 0 0 VDD
port 9 nsew
flabel metal1 2364 1564 2364 1564 0 FreeSans 160 0 0 0 VIP
port 10 nsew
flabel metal1 2380 694 2380 694 0 FreeSans 160 0 0 0 VIN
port 11 nsew
<< end >>
