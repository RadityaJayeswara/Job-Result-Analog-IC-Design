magic
tech sky130A
magscale 1 2
timestamp 1729234290
<< nwell >>
rect 374 -69 1372 2793
<< nsubdiff >>
rect 410 2723 472 2757
rect 1273 2723 1336 2757
rect 410 2697 444 2723
rect 1302 2697 1336 2723
rect 410 1 444 21
rect 1302 1 1336 21
rect 410 -33 472 1
rect 1273 -33 1336 1
<< nsubdiffcont >>
rect 472 2723 1273 2757
rect 410 21 444 2697
rect 1302 21 1336 2697
rect 472 -33 1273 1
<< poly >>
rect 520 2685 586 2701
rect 520 2651 536 2685
rect 570 2651 586 2685
rect 520 2635 586 2651
rect 556 2620 586 2635
rect 1160 2685 1226 2701
rect 1160 2651 1176 2685
rect 1210 2651 1226 2685
rect 1160 2635 1226 2651
rect 1160 2620 1190 2635
rect 520 1989 586 2005
rect 644 2003 844 2109
rect 520 1955 536 1989
rect 570 1955 586 1989
rect 520 1939 586 1955
rect 556 1924 586 1939
rect 1160 1989 1226 2005
rect 1160 1955 1176 1989
rect 1210 1955 1226 1989
rect 1160 1939 1226 1955
rect 1160 1924 1190 1939
rect 644 1310 1102 1412
rect 556 783 586 798
rect 520 767 586 783
rect 520 733 536 767
rect 570 733 586 767
rect 520 717 586 733
rect 1160 783 1190 798
rect 1160 767 1226 783
rect 1160 733 1176 767
rect 1210 733 1226 767
rect 902 614 1102 720
rect 1160 717 1226 733
rect 556 89 586 104
rect 520 73 586 89
rect 520 39 536 73
rect 570 39 586 73
rect 520 23 586 39
rect 1160 89 1190 104
rect 1160 73 1226 89
rect 1160 39 1176 73
rect 1210 39 1226 73
rect 1160 23 1226 39
<< polycont >>
rect 536 2651 570 2685
rect 1176 2651 1210 2685
rect 536 1955 570 1989
rect 1176 1955 1210 1989
rect 536 733 570 767
rect 1176 733 1210 767
rect 536 39 570 73
rect 1176 39 1210 73
<< locali >>
rect 410 2723 472 2757
rect 1273 2723 1336 2757
rect 410 2697 444 2723
rect 1302 2697 1336 2723
rect 520 2651 536 2685
rect 570 2651 586 2685
rect 1160 2651 1176 2685
rect 1210 2651 1226 2685
rect 520 1955 536 1989
rect 570 1955 586 1989
rect 1160 1955 1176 1989
rect 1210 1955 1226 1989
rect 520 733 536 767
rect 570 733 586 767
rect 1160 733 1176 767
rect 1210 733 1226 767
rect 520 39 536 73
rect 570 39 586 73
rect 1160 39 1176 73
rect 1210 39 1226 73
rect 410 1 444 21
rect 1302 1 1336 21
rect 410 -33 472 1
rect 1273 -33 1336 1
<< viali >>
rect 1156 2757 1232 2762
rect 1156 2726 1232 2757
rect 536 2651 570 2685
rect 1176 2651 1210 2685
rect 536 1955 570 1989
rect 1176 1955 1210 1989
rect 536 733 570 767
rect 1176 733 1210 767
rect 536 39 570 73
rect 1176 39 1210 73
rect 510 -33 586 -2
rect 510 -38 586 -33
<< metal1 >>
rect 1144 2762 1244 2768
rect 1144 2726 1156 2762
rect 1232 2726 1244 2762
rect 1144 2720 1244 2726
rect 1164 2691 1236 2720
rect 524 2685 582 2691
rect 1061 2690 1236 2691
rect 524 2684 536 2685
rect 511 2651 536 2684
rect 570 2651 582 2685
rect 511 2645 582 2651
rect 850 2685 1236 2690
rect 850 2651 1176 2685
rect 1210 2651 1236 2685
rect 850 2647 1236 2651
rect 511 2603 545 2645
rect 497 2593 637 2603
rect 491 2216 501 2593
rect 553 2216 637 2593
rect 497 2204 637 2216
rect 524 1989 582 1995
rect 510 1955 536 1989
rect 570 1955 582 1989
rect 510 1949 582 1955
rect 510 1907 544 1949
rect 498 1896 638 1907
rect 498 1520 589 1896
rect 641 1520 651 1896
rect 498 1508 638 1520
rect 592 1255 815 1301
rect 592 1214 638 1255
rect 498 814 638 1214
rect 510 773 544 814
rect 510 767 582 773
rect 510 733 536 767
rect 570 733 582 767
rect 524 727 582 733
rect 498 120 638 520
rect 510 79 544 120
rect 850 79 896 2647
rect 1061 2645 1236 2647
rect 1202 2602 1236 2645
rect 1110 2204 1249 2602
rect 1164 1989 1222 1995
rect 1164 1955 1176 1989
rect 1210 1955 1235 1989
rect 1164 1949 1235 1955
rect 1202 1908 1235 1949
rect 1108 1508 1248 1908
rect 1108 1467 1154 1508
rect 931 1421 1154 1467
rect 1108 1202 1248 1214
rect 1095 826 1105 1202
rect 1157 826 1248 1202
rect 1108 814 1248 826
rect 1202 773 1236 814
rect 1164 767 1236 773
rect 1164 733 1176 767
rect 1210 733 1236 767
rect 1164 727 1222 733
rect 1108 508 1248 520
rect 1108 132 1193 508
rect 1245 132 1255 508
rect 1108 120 1248 132
rect 1203 79 1236 120
rect 510 73 896 79
rect 510 39 536 73
rect 570 39 896 73
rect 510 33 896 39
rect 1164 73 1236 79
rect 1164 39 1176 73
rect 1210 39 1236 73
rect 1164 33 1222 39
rect 510 4 582 33
rect 498 -2 598 4
rect 498 -38 510 -2
rect 586 -38 598 -2
rect 498 -44 598 -38
<< via1 >>
rect 501 2216 553 2593
rect 589 1520 641 1896
rect 1105 826 1157 1202
rect 1193 132 1245 508
<< metal2 >>
rect 501 2593 553 2603
rect 501 2206 553 2216
rect 501 2154 552 2206
rect 504 2093 549 2154
rect 498 2084 554 2093
rect 498 2019 554 2028
rect 1180 2026 1189 2086
rect 1249 2026 1258 2086
rect 504 697 549 2019
rect 589 1896 641 1906
rect 589 1387 641 1520
rect 1105 1387 1157 1388
rect 589 1335 1157 1387
rect 1105 1202 1157 1335
rect 1105 816 1157 826
rect 1193 704 1245 2026
rect 488 637 497 697
rect 557 637 566 697
rect 1192 695 1248 704
rect 1192 630 1248 639
rect 1193 508 1245 630
rect 1193 122 1245 132
<< via2 >>
rect 498 2028 554 2084
rect 1189 2026 1249 2086
rect 497 637 557 697
rect 1192 639 1248 695
<< metal3 >>
rect 493 2086 559 2089
rect 1184 2086 1254 2091
rect 493 2084 1189 2086
rect 493 2028 498 2084
rect 554 2028 1189 2084
rect 493 2026 1189 2028
rect 1249 2026 1254 2086
rect 493 2023 559 2026
rect 1184 2021 1254 2026
rect 492 697 562 702
rect 1187 697 1253 700
rect 492 637 497 697
rect 557 695 1253 697
rect 557 639 1192 695
rect 1248 639 1253 695
rect 557 637 1253 639
rect 492 632 562 637
rect 1187 634 1253 637
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729132701
transform 1 0 571 0 1 1014
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729132701
transform 1 0 1175 0 1 2404
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729132701
transform 1 0 1175 0 1 1708
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729132701
transform 1 0 1175 0 1 1014
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729132701
transform 1 0 1175 0 1 320
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729132701
transform 1 0 571 0 1 320
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729132701
transform 1 0 571 0 1 1708
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729132701
transform 1 0 571 0 1 2404
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729141730
transform 1 0 873 0 1 2404
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729141730
transform 1 0 873 0 1 1708
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729141730
transform 1 0 873 0 1 1014
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729141730
transform 1 0 873 0 1 320
box -323 -300 323 300
<< labels >>
flabel metal1 1178 2474 1178 2474 0 FreeSans 240 0 0 0 VDD
port 2 nsew
flabel metal1 574 930 574 930 0 FreeSans 240 0 0 0 D2
port 4 nsew
flabel metal2 1226 710 1226 710 0 FreeSans 240 0 0 0 D5
port 7 nsew
flabel metal2 612 1472 612 1472 0 FreeSans 240 0 0 0 D1
port 8 nsew
<< end >>
