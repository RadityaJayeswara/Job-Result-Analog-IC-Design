magic
tech sky130A
magscale 1 2
timestamp 1729223995
<< nmos >>
rect -407 109 -247 309
rect -189 109 -29 309
rect 29 109 189 309
rect 247 109 407 309
rect -407 -309 -247 -109
rect -189 -309 -29 -109
rect 29 -309 189 -109
rect 247 -309 407 -109
<< ndiff >>
rect -465 297 -407 309
rect -465 121 -453 297
rect -419 121 -407 297
rect -465 109 -407 121
rect -247 297 -189 309
rect -247 121 -235 297
rect -201 121 -189 297
rect -247 109 -189 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 189 297 247 309
rect 189 121 201 297
rect 235 121 247 297
rect 189 109 247 121
rect 407 297 465 309
rect 407 121 419 297
rect 453 121 465 297
rect 407 109 465 121
rect -465 -121 -407 -109
rect -465 -297 -453 -121
rect -419 -297 -407 -121
rect -465 -309 -407 -297
rect -247 -121 -189 -109
rect -247 -297 -235 -121
rect -201 -297 -189 -121
rect -247 -309 -189 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 189 -121 247 -109
rect 189 -297 201 -121
rect 235 -297 247 -121
rect 189 -309 247 -297
rect 407 -121 465 -109
rect 407 -297 419 -121
rect 453 -297 465 -121
rect 407 -309 465 -297
<< ndiffc >>
rect -453 121 -419 297
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect 419 121 453 297
rect -453 -297 -419 -121
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect 419 -297 453 -121
<< poly >>
rect -407 381 -247 397
rect -407 347 -391 381
rect -263 347 -247 381
rect -407 309 -247 347
rect -189 381 -29 397
rect -189 347 -173 381
rect -45 347 -29 381
rect -189 309 -29 347
rect 29 381 189 397
rect 29 347 45 381
rect 173 347 189 381
rect 29 309 189 347
rect 247 381 407 397
rect 247 347 263 381
rect 391 347 407 381
rect 247 309 407 347
rect -407 71 -247 109
rect -407 37 -391 71
rect -263 37 -247 71
rect -407 21 -247 37
rect -189 71 -29 109
rect -189 37 -173 71
rect -45 37 -29 71
rect -189 21 -29 37
rect 29 71 189 109
rect 29 37 45 71
rect 173 37 189 71
rect 29 21 189 37
rect 247 71 407 109
rect 247 37 263 71
rect 391 37 407 71
rect 247 21 407 37
rect -407 -37 -247 -21
rect -407 -71 -391 -37
rect -263 -71 -247 -37
rect -407 -109 -247 -71
rect -189 -37 -29 -21
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect -189 -109 -29 -71
rect 29 -37 189 -21
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 29 -109 189 -71
rect 247 -37 407 -21
rect 247 -71 263 -37
rect 391 -71 407 -37
rect 247 -109 407 -71
rect -407 -347 -247 -309
rect -407 -381 -391 -347
rect -263 -381 -247 -347
rect -407 -397 -247 -381
rect -189 -347 -29 -309
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect -189 -397 -29 -381
rect 29 -347 189 -309
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 29 -397 189 -381
rect 247 -347 407 -309
rect 247 -381 263 -347
rect 391 -381 407 -347
rect 247 -397 407 -381
<< polycont >>
rect -391 347 -263 381
rect -173 347 -45 381
rect 45 347 173 381
rect 263 347 391 381
rect -391 37 -263 71
rect -173 37 -45 71
rect 45 37 173 71
rect 263 37 391 71
rect -391 -71 -263 -37
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect 263 -71 391 -37
rect -391 -381 -263 -347
rect -173 -381 -45 -347
rect 45 -381 173 -347
rect 263 -381 391 -347
<< locali >>
rect -407 347 -391 381
rect -263 347 -247 381
rect -189 347 -173 381
rect -45 347 -29 381
rect 29 347 45 381
rect 173 347 189 381
rect 247 347 263 381
rect 391 347 407 381
rect -453 297 -419 313
rect -453 105 -419 121
rect -235 297 -201 313
rect -235 105 -201 121
rect -17 297 17 313
rect -17 105 17 121
rect 201 297 235 313
rect 201 105 235 121
rect 419 297 453 313
rect 419 105 453 121
rect -407 37 -391 71
rect -263 37 -247 71
rect -189 37 -173 71
rect -45 37 -29 71
rect 29 37 45 71
rect 173 37 189 71
rect 247 37 263 71
rect 391 37 407 71
rect -407 -71 -391 -37
rect -263 -71 -247 -37
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 247 -71 263 -37
rect 391 -71 407 -37
rect -453 -121 -419 -105
rect -453 -313 -419 -297
rect -235 -121 -201 -105
rect -235 -313 -201 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 201 -121 235 -105
rect 201 -313 235 -297
rect 419 -121 453 -105
rect 419 -313 453 -297
rect -407 -381 -391 -347
rect -263 -381 -247 -347
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 247 -381 263 -347
rect 391 -381 407 -347
<< viali >>
rect -391 347 -263 381
rect -173 347 -45 381
rect 45 347 173 381
rect 263 347 391 381
rect -453 121 -419 297
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect 419 121 453 297
rect -391 37 -263 71
rect -173 37 -45 71
rect 45 37 173 71
rect 263 37 391 71
rect -391 -71 -263 -37
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect 263 -71 391 -37
rect -453 -297 -419 -121
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect 419 -297 453 -121
rect -391 -381 -263 -347
rect -173 -381 -45 -347
rect 45 -381 173 -347
rect 263 -381 391 -347
<< metal1 >>
rect -403 381 -251 387
rect -403 347 -391 381
rect -263 347 -251 381
rect -403 341 -251 347
rect -185 381 -33 387
rect -185 347 -173 381
rect -45 347 -33 381
rect -185 341 -33 347
rect 33 381 185 387
rect 33 347 45 381
rect 173 347 185 381
rect 33 341 185 347
rect 251 381 403 387
rect 251 347 263 381
rect 391 347 403 381
rect 251 341 403 347
rect -459 297 -413 309
rect -459 121 -453 297
rect -419 121 -413 297
rect -459 109 -413 121
rect -241 297 -195 309
rect -241 121 -235 297
rect -201 121 -195 297
rect -241 109 -195 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 195 297 241 309
rect 195 121 201 297
rect 235 121 241 297
rect 195 109 241 121
rect 413 297 459 309
rect 413 121 419 297
rect 453 121 459 297
rect 413 109 459 121
rect -403 71 -251 77
rect -403 37 -391 71
rect -263 37 -251 71
rect -403 31 -251 37
rect -185 71 -33 77
rect -185 37 -173 71
rect -45 37 -33 71
rect -185 31 -33 37
rect 33 71 185 77
rect 33 37 45 71
rect 173 37 185 71
rect 33 31 185 37
rect 251 71 403 77
rect 251 37 263 71
rect 391 37 403 71
rect 251 31 403 37
rect -403 -37 -251 -31
rect -403 -71 -391 -37
rect -263 -71 -251 -37
rect -403 -77 -251 -71
rect -185 -37 -33 -31
rect -185 -71 -173 -37
rect -45 -71 -33 -37
rect -185 -77 -33 -71
rect 33 -37 185 -31
rect 33 -71 45 -37
rect 173 -71 185 -37
rect 33 -77 185 -71
rect 251 -37 403 -31
rect 251 -71 263 -37
rect 391 -71 403 -37
rect 251 -77 403 -71
rect -459 -121 -413 -109
rect -459 -297 -453 -121
rect -419 -297 -413 -121
rect -459 -309 -413 -297
rect -241 -121 -195 -109
rect -241 -297 -235 -121
rect -201 -297 -195 -121
rect -241 -309 -195 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 195 -121 241 -109
rect 195 -297 201 -121
rect 235 -297 241 -121
rect 195 -309 241 -297
rect 413 -121 459 -109
rect 413 -297 419 -121
rect 453 -297 459 -121
rect 413 -309 459 -297
rect -403 -347 -251 -341
rect -403 -381 -391 -347
rect -263 -381 -251 -347
rect -403 -387 -251 -381
rect -185 -347 -33 -341
rect -185 -381 -173 -347
rect -45 -381 -33 -347
rect -185 -387 -33 -381
rect 33 -347 185 -341
rect 33 -381 45 -347
rect 173 -381 185 -347
rect 33 -387 185 -381
rect 251 -347 403 -341
rect 251 -381 263 -347
rect 391 -381 403 -347
rect 251 -387 403 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
