magic
tech sky130A
magscale 1 2
timestamp 1729410161
<< nwell >>
rect -4586 1118 -3594 1866
<< viali >>
rect -3660 644 -3626 726
rect -3558 644 -3524 726
rect -3422 404 -3283 527
rect -3420 196 -3281 320
rect -3421 -27 -3282 97
rect -3660 -214 -3626 -147
rect -3421 -242 -3282 -118
rect -3419 -426 -3280 -302
rect -3420 -660 -3281 -536
rect -3136 -632 -3102 -564
<< metal1 >>
rect -4437 1210 -2977 1267
rect -4437 970 -4380 1210
rect -3666 726 -3518 738
rect -3666 644 -3660 726
rect -3626 644 -3558 726
rect -3524 644 -3518 726
rect -3666 632 -3518 644
rect -3382 533 -3324 897
rect -3434 527 -3271 533
rect -3434 404 -3422 527
rect -3283 404 -3271 527
rect -3434 398 -3271 404
rect -3432 320 -3269 326
rect -3432 196 -3420 320
rect -3281 196 -3269 320
rect -3432 190 -3269 196
rect -3433 97 -3270 103
rect -3433 -27 -3421 97
rect -3282 69 -3270 97
rect -3178 69 -3110 814
rect -2158 642 -2112 921
rect -2494 596 -2112 642
rect -2494 383 -2448 596
rect -3031 195 -3021 371
rect -2969 195 -2959 371
rect -3282 1 -3110 69
rect -3282 -27 -3270 1
rect -3433 -33 -3270 -27
rect -3433 -118 -3270 -112
rect -3433 -135 -3421 -118
rect -3666 -147 -3421 -135
rect -3666 -214 -3660 -147
rect -3626 -214 -3421 -147
rect -3666 -226 -3421 -214
rect -3433 -242 -3421 -226
rect -3282 -242 -3270 -118
rect -3433 -248 -3270 -242
rect -3431 -302 -3268 -296
rect -3431 -426 -3419 -302
rect -3280 -426 -3268 -302
rect -2718 -356 -2512 -286
rect -3431 -432 -3268 -426
rect -3432 -536 -3269 -529
rect -3432 -660 -3420 -536
rect -3281 -552 -3269 -536
rect -3281 -564 -3096 -552
rect -3281 -632 -3136 -564
rect -3102 -632 -3096 -564
rect -3281 -644 -3096 -632
rect -3281 -660 -3269 -644
rect -3432 -666 -3269 -660
rect -3714 -763 -3048 -704
rect -4031 -978 -3889 -948
rect -4031 -979 -3860 -978
rect -4031 -1038 -2990 -979
rect -4031 -1068 -3889 -1038
rect -3049 -1191 -2990 -1038
<< via1 >>
rect -3420 196 -3281 320
rect -3021 195 -2969 371
rect -3419 -426 -3280 -302
<< metal2 >>
rect -2740 1083 -2684 1093
rect -2740 897 -2684 907
rect -3420 320 -3281 330
rect -3182 295 -3110 695
rect -3281 223 -3110 295
rect -3023 371 -2967 381
rect -3420 186 -3281 196
rect -3023 185 -2967 195
rect -3419 -302 -3280 -292
rect -3280 -394 -2393 -342
rect -3419 -436 -3280 -426
rect -2445 -517 -2393 -394
rect -2444 -530 -2393 -517
<< via2 >>
rect -2740 907 -2684 1083
rect -3023 195 -3021 371
rect -3021 195 -2969 371
rect -2969 195 -2967 371
<< metal3 >>
rect -2750 1083 -2674 1088
rect -2750 907 -2740 1083
rect -2684 907 -2674 1083
rect -2750 629 -2674 907
rect -3033 553 -2674 629
rect -3033 371 -2957 553
rect -3033 195 -3023 371
rect -2967 195 -2957 371
rect -3033 190 -2957 195
use biasdif  biasdif_0
timestamp 1729225851
transform 1 0 -3263 0 1 -842
box 151 556 1433 1384
use difpair  difpair_0
timestamp 1729394227
transform 1 0 -5088 0 1 99
box 1494 509 3258 1768
use nmoscsi  nmoscsi_0
timestamp 1729218094
transform 1 0 -2834 0 1 -1003
box -302 -747 1004 647
use pmoscs  pmoscs_0
timestamp 1729234290
transform 1 0 -4962 0 1 -1675
box 374 -69 1372 2793
<< labels >>
flabel metal1 -3205 -740 -3205 -740 0 FreeSans 640 0 0 0 D1-3
flabel metal1 -3181 -1005 -3181 -1005 0 FreeSans 640 0 0 0 D2-4
flabel space -2777 593 -2777 593 0 FreeSans 640 0 0 0 D6-8-M9
flabel metal1 -2133 620 -2133 620 0 FreeSans 640 0 0 0 D7-9
flabel viali -3352 463 -3352 463 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel via1 -3351 255 -3351 255 0 FreeSans 640 0 0 0 VIN
port 2 nsew
flabel viali -3355 31 -3355 31 0 FreeSans 640 0 0 0 VIP
port 3 nsew
flabel viali -3348 -185 -3348 -185 0 FreeSans 640 0 0 0 VDD
port 4 nsew
flabel viali -3345 -363 -3345 -363 0 FreeSans 640 0 0 0 RS
port 5 nsew
flabel viali -3352 -600 -3352 -600 0 FreeSans 640 0 0 0 GND
port 7 nsew
<< end >>
