magic
tech sky130A
magscale 1 2
timestamp 1729135101
<< nwell >>
rect -323 -300 323 300
<< pmos >>
rect -229 -200 -29 200
rect 29 -200 229 200
<< pdiff >>
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
<< pdiffc >>
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
<< poly >>
rect -208 281 -50 297
rect -208 264 -192 281
rect -229 247 -192 264
rect -66 264 -50 281
rect 50 281 208 297
rect 50 264 66 281
rect -66 247 -29 264
rect -229 200 -29 247
rect 29 247 66 264
rect 192 264 208 281
rect 192 247 229 264
rect 29 200 229 247
rect -229 -247 -29 -200
rect -229 -264 -192 -247
rect -208 -281 -192 -264
rect -66 -264 -29 -247
rect 29 -247 229 -200
rect 29 -264 66 -247
rect -66 -281 -50 -264
rect -208 -297 -50 -281
rect 50 -281 66 -264
rect 192 -264 229 -247
rect 192 -281 208 -264
rect 50 -297 208 -281
<< polycont >>
rect -192 247 -66 281
rect 66 247 192 281
rect -192 -281 -66 -247
rect 66 -281 192 -247
<< locali >>
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
<< viali >>
rect -213 247 -192 281
rect -192 247 -66 281
rect -66 247 -45 281
rect 45 247 66 281
rect 66 247 192 281
rect 192 247 213 281
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect -213 -281 -192 -247
rect -192 -281 -66 -247
rect -66 -281 -45 -247
rect 45 -281 66 -247
rect 66 -281 192 -247
rect 192 -281 213 -247
<< metal1 >>
rect -225 281 -33 287
rect -225 247 -213 281
rect -45 247 -33 281
rect -225 241 -33 247
rect 33 281 225 287
rect 33 247 45 281
rect 213 247 225 281
rect 33 241 225 247
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect -225 -247 -33 -241
rect -225 -281 -213 -247
rect -45 -281 -33 -247
rect -225 -287 -33 -281
rect 33 -247 225 -241
rect 33 -281 45 -247
rect 213 -281 225 -247
rect 33 -287 225 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 75 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
