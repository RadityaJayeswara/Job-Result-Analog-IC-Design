magic
tech sky130A
magscale 1 2
timestamp 1729233515
<< error_p >>
rect -223 454 223 672
rect -223 18 223 236
rect -223 -418 223 -200
<< nwell >>
rect -223 454 223 854
rect -223 18 223 418
rect -223 -418 223 -18
rect -223 -854 223 -454
<< pmos >>
rect -129 554 -29 754
rect 29 554 129 754
rect -129 118 -29 318
rect 29 118 129 318
rect -129 -318 -29 -118
rect 29 -318 129 -118
rect -129 -754 -29 -554
rect 29 -754 129 -554
<< pdiff >>
rect -187 742 -129 754
rect -187 566 -175 742
rect -141 566 -129 742
rect -187 554 -129 566
rect -29 742 29 754
rect -29 566 -17 742
rect 17 566 29 742
rect -29 554 29 566
rect 129 742 187 754
rect 129 566 141 742
rect 175 566 187 742
rect 129 554 187 566
rect -187 306 -129 318
rect -187 130 -175 306
rect -141 130 -129 306
rect -187 118 -129 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 129 306 187 318
rect 129 130 141 306
rect 175 130 187 306
rect 129 118 187 130
rect -187 -130 -129 -118
rect -187 -306 -175 -130
rect -141 -306 -129 -130
rect -187 -318 -129 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 129 -130 187 -118
rect 129 -306 141 -130
rect 175 -306 187 -130
rect 129 -318 187 -306
rect -187 -566 -129 -554
rect -187 -742 -175 -566
rect -141 -742 -129 -566
rect -187 -754 -129 -742
rect -29 -566 29 -554
rect -29 -742 -17 -566
rect 17 -742 29 -566
rect -29 -754 29 -742
rect 129 -566 187 -554
rect 129 -742 141 -566
rect 175 -742 187 -566
rect 129 -754 187 -742
<< pdiffc >>
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
<< poly >>
rect -129 835 -29 851
rect -129 801 -113 835
rect -45 801 -29 835
rect -129 754 -29 801
rect 29 835 129 851
rect 29 801 45 835
rect 113 801 129 835
rect 29 754 129 801
rect -129 507 -29 554
rect -129 473 -113 507
rect -45 473 -29 507
rect -129 457 -29 473
rect 29 507 129 554
rect 29 473 45 507
rect 113 473 129 507
rect 29 457 129 473
rect -129 399 -29 415
rect -129 365 -113 399
rect -45 365 -29 399
rect -129 318 -29 365
rect 29 399 129 415
rect 29 365 45 399
rect 113 365 129 399
rect 29 318 129 365
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect -129 -365 -29 -318
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect -129 -415 -29 -399
rect 29 -365 129 -318
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 29 -415 129 -399
rect -129 -473 -29 -457
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect -129 -554 -29 -507
rect 29 -473 129 -457
rect 29 -507 45 -473
rect 113 -507 129 -473
rect 29 -554 129 -507
rect -129 -801 -29 -754
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect -129 -851 -29 -835
rect 29 -801 129 -754
rect 29 -835 45 -801
rect 113 -835 129 -801
rect 29 -851 129 -835
<< polycont >>
rect -113 801 -45 835
rect 45 801 113 835
rect -113 473 -45 507
rect 45 473 113 507
rect -113 365 -45 399
rect 45 365 113 399
rect -113 37 -45 71
rect 45 37 113 71
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect -113 -507 -45 -473
rect 45 -507 113 -473
rect -113 -835 -45 -801
rect 45 -835 113 -801
<< locali >>
rect -129 801 -113 835
rect -45 801 -29 835
rect 29 801 45 835
rect 113 801 129 835
rect -175 742 -141 758
rect -175 550 -141 566
rect -17 742 17 758
rect -17 550 17 566
rect 141 742 175 758
rect 141 550 175 566
rect -129 473 -113 507
rect -45 473 -29 507
rect 29 473 45 507
rect 113 473 129 507
rect -129 365 -113 399
rect -45 365 -29 399
rect 29 365 45 399
rect 113 365 129 399
rect -175 306 -141 322
rect -175 114 -141 130
rect -17 306 17 322
rect -17 114 17 130
rect 141 306 175 322
rect 141 114 175 130
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect -175 -130 -141 -114
rect -175 -322 -141 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 141 -130 175 -114
rect 141 -322 175 -306
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 113 -399 129 -365
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect 29 -507 45 -473
rect 113 -507 129 -473
rect -175 -566 -141 -550
rect -175 -758 -141 -742
rect -17 -566 17 -550
rect -17 -758 17 -742
rect 141 -566 175 -550
rect 141 -758 175 -742
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect 29 -835 45 -801
rect 113 -835 129 -801
<< viali >>
rect -105 801 -53 835
rect 53 801 105 835
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect -105 473 -53 507
rect 53 473 105 507
rect -105 365 -53 399
rect 53 365 105 399
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect -105 37 -53 71
rect 53 37 105 71
rect -105 -71 -53 -37
rect 53 -71 105 -37
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect -105 -399 -53 -365
rect 53 -399 105 -365
rect -105 -507 -53 -473
rect 53 -507 105 -473
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
rect -105 -835 -53 -801
rect 53 -835 105 -801
<< metal1 >>
rect -117 835 -41 841
rect -117 801 -105 835
rect -53 801 -41 835
rect -117 795 -41 801
rect 41 835 117 841
rect 41 801 53 835
rect 105 801 117 835
rect 41 795 117 801
rect -181 742 -135 754
rect -181 566 -175 742
rect -141 566 -135 742
rect -181 554 -135 566
rect -23 742 23 754
rect -23 566 -17 742
rect 17 566 23 742
rect -23 554 23 566
rect 135 742 181 754
rect 135 566 141 742
rect 175 566 181 742
rect 135 554 181 566
rect -117 507 -41 513
rect -117 473 -105 507
rect -53 473 -41 507
rect -117 467 -41 473
rect 41 507 117 513
rect 41 473 53 507
rect 105 473 117 507
rect 41 467 117 473
rect -117 399 -41 405
rect -117 365 -105 399
rect -53 365 -41 399
rect -117 359 -41 365
rect 41 399 117 405
rect 41 365 53 399
rect 105 365 117 399
rect 41 359 117 365
rect -181 306 -135 318
rect -181 130 -175 306
rect -141 130 -135 306
rect -181 118 -135 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 135 306 181 318
rect 135 130 141 306
rect 175 130 181 306
rect 135 118 181 130
rect -117 71 -41 77
rect -117 37 -105 71
rect -53 37 -41 71
rect -117 31 -41 37
rect 41 71 117 77
rect 41 37 53 71
rect 105 37 117 71
rect 41 31 117 37
rect -117 -37 -41 -31
rect -117 -71 -105 -37
rect -53 -71 -41 -37
rect -117 -77 -41 -71
rect 41 -37 117 -31
rect 41 -71 53 -37
rect 105 -71 117 -37
rect 41 -77 117 -71
rect -181 -130 -135 -118
rect -181 -306 -175 -130
rect -141 -306 -135 -130
rect -181 -318 -135 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 135 -130 181 -118
rect 135 -306 141 -130
rect 175 -306 181 -130
rect 135 -318 181 -306
rect -117 -365 -41 -359
rect -117 -399 -105 -365
rect -53 -399 -41 -365
rect -117 -405 -41 -399
rect 41 -365 117 -359
rect 41 -399 53 -365
rect 105 -399 117 -365
rect 41 -405 117 -399
rect -117 -473 -41 -467
rect -117 -507 -105 -473
rect -53 -507 -41 -473
rect -117 -513 -41 -507
rect 41 -473 117 -467
rect 41 -507 53 -473
rect 105 -507 117 -473
rect 41 -513 117 -507
rect -181 -566 -135 -554
rect -181 -742 -175 -566
rect -141 -742 -135 -566
rect -181 -754 -135 -742
rect -23 -566 23 -554
rect -23 -742 -17 -566
rect 17 -742 23 -566
rect -23 -754 23 -742
rect 135 -566 181 -554
rect 135 -742 141 -566
rect 175 -742 181 -566
rect 135 -754 181 -742
rect -117 -801 -41 -795
rect -117 -835 -105 -801
rect -53 -835 -41 -801
rect -117 -841 -41 -835
rect 41 -801 117 -795
rect 41 -835 53 -801
rect 105 -835 117 -801
rect 41 -841 117 -835
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
