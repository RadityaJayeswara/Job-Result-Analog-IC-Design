magic
tech sky130A
magscale 1 2
timestamp 1728978902
<< error_p >>
rect -29 -61 29 -55
rect -29 -95 -17 -61
rect -29 -101 29 -95
<< nwell >>
rect -211 -234 211 234
<< pmos >>
rect -15 -14 15 86
<< pdiff >>
rect -73 74 -15 86
rect -73 -2 -61 74
rect -27 -2 -15 74
rect -73 -14 -15 -2
rect 15 74 73 86
rect 15 -2 27 74
rect 61 -2 73 74
rect 15 -14 73 -2
<< pdiffc >>
rect -61 -2 -27 74
rect 27 -2 61 74
<< nsubdiff >>
rect -175 164 -79 198
rect 79 164 175 198
rect -175 101 -141 164
rect 141 101 175 164
rect -175 -164 -141 -101
rect 141 -164 175 -101
rect -175 -198 -79 -164
rect 79 -198 175 -164
<< nsubdiffcont >>
rect -79 164 79 198
rect -175 -101 -141 101
rect 141 -101 175 101
rect -79 -198 79 -164
<< poly >>
rect -15 86 15 112
rect -15 -45 15 -14
rect -33 -61 33 -45
rect -33 -95 -17 -61
rect 17 -95 33 -61
rect -33 -111 33 -95
<< polycont >>
rect -17 -95 17 -61
<< locali >>
rect -175 164 -79 198
rect 79 164 175 198
rect -175 101 -141 164
rect 141 101 175 164
rect -61 74 -27 90
rect -61 -18 -27 -2
rect 27 74 61 90
rect 27 -18 61 -2
rect -33 -95 -17 -61
rect 17 -95 33 -61
rect -175 -164 -141 -101
rect 141 -164 175 -101
rect -175 -198 -79 -164
rect 79 -198 175 -164
<< viali >>
rect -61 -2 -27 74
rect 27 -2 61 74
rect -17 -95 17 -61
<< metal1 >>
rect -67 74 -21 86
rect -67 -2 -61 74
rect -27 -2 -21 74
rect -67 -14 -21 -2
rect 21 74 67 86
rect 21 -2 27 74
rect 61 -2 67 74
rect 21 -14 67 -2
rect -29 -61 29 -55
rect -29 -95 -17 -61
rect 17 -95 29 -61
rect -29 -101 29 -95
<< properties >>
string FIXED_BBOX -158 -181 158 181
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
