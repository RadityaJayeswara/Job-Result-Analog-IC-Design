magic
tech sky130A
magscale 1 2
timestamp 1729225851
<< psubdiff >>
rect 151 1344 211 1378
rect 1373 1344 1433 1378
rect 151 1318 185 1344
rect 1399 1318 1433 1344
rect 151 596 185 622
rect 1399 596 1433 622
rect 151 562 211 596
rect 1373 562 1433 596
<< psubdiffcont >>
rect 211 1344 1373 1378
rect 151 622 185 1318
rect 1399 622 1433 1318
rect 211 562 1373 596
<< poly >>
rect 235 1297 327 1313
rect 235 1263 251 1297
rect 285 1263 327 1297
rect 235 1247 327 1263
rect 1257 1297 1349 1313
rect 1257 1263 1299 1297
rect 1333 1263 1349 1297
rect 1257 1247 1349 1263
rect 1257 1225 1287 1247
rect 235 677 327 693
rect 235 643 251 677
rect 285 643 327 677
rect 235 627 327 643
rect 1257 677 1349 693
rect 1257 643 1299 677
rect 1333 643 1349 677
rect 1257 627 1349 643
<< polycont >>
rect 251 1263 285 1297
rect 1299 1263 1333 1297
rect 251 643 285 677
rect 1299 643 1333 677
<< locali >>
rect 151 1344 211 1378
rect 1373 1344 1433 1378
rect 151 1318 185 1344
rect 1399 1318 1433 1344
rect 235 1263 251 1297
rect 285 1263 301 1297
rect 1283 1263 1299 1297
rect 1333 1263 1349 1297
rect 235 643 251 677
rect 285 643 301 677
rect 1283 643 1299 677
rect 1333 643 1349 677
rect 151 596 185 622
rect 1399 596 1433 622
rect 151 562 211 596
rect 1373 562 1433 596
<< viali >>
rect 557 1344 591 1378
rect 993 1344 1027 1378
rect 251 1263 285 1297
rect 1299 1263 1333 1297
rect 251 643 285 677
rect 1299 643 1333 677
rect 557 562 591 596
rect 993 562 1027 596
<< metal1 >>
rect 545 1378 603 1384
rect 545 1344 557 1378
rect 591 1344 603 1378
rect 545 1338 603 1344
rect 981 1378 1039 1384
rect 981 1344 993 1378
rect 1027 1344 1039 1378
rect 981 1338 1039 1344
rect 239 1297 297 1303
rect 239 1263 251 1297
rect 285 1263 297 1297
rect 239 1257 297 1263
rect 245 1225 291 1257
rect 551 1225 597 1338
rect 987 1225 1033 1338
rect 1287 1297 1345 1303
rect 1287 1263 1299 1297
rect 1333 1263 1345 1297
rect 1287 1257 1345 1263
rect 1293 1225 1339 1257
rect 239 1025 379 1225
rect 756 1037 766 1213
rect 818 1037 828 1213
rect 333 993 379 1025
rect 1205 1025 1345 1225
rect 1205 993 1251 1025
rect 333 947 1251 993
rect 769 915 815 947
rect 239 903 379 915
rect 1205 903 1345 915
rect 239 727 330 903
rect 382 727 392 903
rect 1192 727 1202 903
rect 1254 727 1345 903
rect 239 715 379 727
rect 1205 715 1345 727
rect 245 683 291 715
rect 239 677 297 683
rect 239 643 251 677
rect 285 643 297 677
rect 239 637 297 643
rect 551 602 597 715
rect 987 602 1033 715
rect 1293 683 1339 715
rect 1287 677 1345 683
rect 1287 643 1299 677
rect 1333 643 1345 677
rect 1287 637 1345 643
rect 545 596 603 602
rect 545 562 557 596
rect 591 562 603 596
rect 545 556 603 562
rect 981 596 1039 602
rect 981 562 993 596
rect 1027 562 1039 596
rect 981 556 1039 562
<< via1 >>
rect 766 1037 818 1213
rect 330 727 382 903
rect 1202 727 1254 903
<< metal2 >>
rect 766 1213 818 1223
rect 766 996 818 1037
rect 330 944 1254 996
rect 330 903 382 944
rect 330 717 382 727
rect 1202 903 1254 944
rect 1202 717 1254 727
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729223995
transform 1 0 1272 0 1 815
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729223995
transform 1 0 312 0 1 1125
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729223995
transform 1 0 312 0 1 815
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729223995
transform 1 0 1272 0 1 1125
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_YYNGNX  sky130_fd_pr__nfet_01v8_YYNGNX_0
timestamp 1729225706
transform 1 0 792 0 1 970
box -465 -343 465 343
<< labels >>
flabel space 460 1134 460 1134 0 FreeSans 160 0 0 0 M8
flabel space 1116 1132 1116 1132 0 FreeSans 160 0 0 0 M8
flabel space 450 788 450 788 0 FreeSans 160 0 0 0 M9
flabel space 1116 802 1116 802 0 FreeSans 160 0 0 0 M9
flabel space 692 1118 692 1118 0 FreeSans 160 0 0 0 M9
flabel space 904 1120 904 1120 0 FreeSans 160 0 0 0 M9
flabel space 680 810 680 810 0 FreeSans 160 0 0 0 M8
flabel space 900 810 900 810 0 FreeSans 160 0 0 0 M8
flabel via1 793 1125 793 1125 0 FreeSans 160 0 0 0 d9
flabel space 794 811 794 811 0 FreeSans 160 0 0 0 d8
flabel via1 359 811 359 811 0 FreeSans 160 0 0 0 d9
flabel space 575 816 575 816 0 FreeSans 160 0 0 0 S
flabel space 575 1127 575 1127 0 FreeSans 160 0 0 0 S
flabel space 1008 1126 1008 1126 0 FreeSans 160 0 0 0 S
flabel space 1010 813 1010 813 0 FreeSans 160 0 0 0 S
flabel metal1 573 1309 573 1309 0 FreeSans 160 0 0 0 GND
port 1 nsew
flabel metal2 1226 928 1226 928 0 FreeSans 160 0 0 0 D9
port 2 nsew
flabel metal1 1228 1011 1228 1011 0 FreeSans 160 0 0 0 D8
port 3 nsew
<< end >>
